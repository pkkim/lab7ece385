//HDMI Text Controller Example Testbench for ECE 385
//Spring 2024 Distribution

//Modified 3/10/24 by Zuofu
//
//Based on Realdigital documentation on simulating AXI Bus
//as well as BMP writing code from @BrianHGinc
//
//Used for simulation of AXI4-Lite bus as well as generating
//simulation video image for testing

`define SIM_VIDEO //Comment out to simulate AXI bus only
                    //Uncomment to simulate entire screen and write BMP (slow)

module hdmi_text_controller_tb();

	//clock and reset_n signals
	logic aclk =1'b0;
	logic arstn = 1'b0;
	
	//Write Address channel (AW)
	logic [31:0] write_addr =32'd0;	//Master write address
	logic [2:0] write_prot = 3'd0;	//type of write(leave at 0)
	logic write_addr_valid = 1'b0;	//master indicating address is valid
	logic write_addr_ready;		    //slave ready to receive address

	//Write Data Channel (W)
	logic [31:0] write_data = 32'd0;	//Master write data
	logic [3:0] write_strb = 4'd0;	    //Master byte-wise write strobe
	logic write_data_valid = 1'b0;	    //Master indicating write data is valid
	logic write_data_ready;		        //slave ready to receive data

	//Write Response Channel (WR)
	logic write_resp_ready = 1'b0;	//Master ready to receive write response
	logic [1:0] write_resp;		    //slave write response
	logic write_resp_valid;		    //slave response valid
	
	//Read Address channel (AR)
	logic [31:0] read_addr = 32'd0;	//Master read address
	logic [2:0] read_prot =3'd0;	//type of read(leave at 0)
	logic read_addr_valid = 1'b0;	//Master indicating address is valid
	logic read_addr_ready;		    //slave ready to receive address

	//Read Data Channel (R)
	logic read_data_ready = 1'b0;	//Master indicating ready to receive data
	logic [31:0] read_data;		    //slave read data
	logic [1:0] read_resp;		    //slave read response
	logic read_data_valid;		    //slave indicating data in channel is valid

    //Although we can look at the HDMI signal, it is not particularly useful for debugging
    //Instead, simulate and record the pixel clock and the pixel RGB values to generate
    //a simulated image
    logic [3:0] pixel_rgb [3];
    logic pixel_clk, pixel_hs, pixel_vs, pixel_vde;
    logic [9:0] drawX, drawY;
    logic [31:0] tb_read;
    
    //BMP writer related signals    
    localparam BMP_WIDTH  = 800;
    localparam BMP_HEIGHT = 525;
    logic [23:0] bitmap [BMP_WIDTH][BMP_HEIGHT];

    integer i,j; //use integers for loop indices, etc

	//Instantiation of DUT (HDMI TEXT_CONTROLLER) IP
	hdmi_text_controller_v1_0 # (
		.C_AXI_DATA_WIDTH(32),
		.C_AXI_ADDR_WIDTH(16)
	) hdmi_text_controller_v1_0_inst (

		.axi_aclk(aclk),
		.axi_aresetn(arstn),

		.axi_awaddr(write_addr),
		.axi_awprot(write_prot),
		.axi_awvalid(write_addr_valid),
		.axi_awready(write_addr_ready),

		.axi_wdata(write_data),
		.axi_wstrb(write_strb),
		.axi_wvalid(write_data_valid),
		.axi_wready(write_data_ready),

		.axi_bresp(write_resp),
		.axi_bvalid(write_resp_valid),
		.axi_bready(write_resp_ready),

		.axi_araddr(read_addr),
		.axi_arprot(read_prot),
		.axi_arvalid(read_addr_valid),
		.axi_arready(read_addr_ready),

		.axi_rdata(read_data),
		.axi_rresp(read_resp),
		.axi_rvalid(read_data_valid),
		.axi_rready(read_data_ready)
	);
	
	initial begin: CLOCK_INITIALIZATION
	   aclk = 1'b1;
    end 
       
    always begin : CLOCK_GENERATION
        #5 aclk = ~aclk;
    end

    //Uncomment and fill in the following with your own hierarchical reference (e.g. internal signals) 
    //so that the testbench can properly reflect the pixels being draw. 
    //Note that looking at the HDMI signal is not particularly useful here, as it is difficult
    //to decode. E.g. if your hdmi_text_controller has an internal signal named 'clk_25MHz' for
    //the pixel clock, assign pixel_clk = hdmi_text_controller_v1_0_inst.clk_25MHz
    
    // Red Green and Blue values respectively - these come from your draw logic
     assign pixel_rgb[0] = hdmi_text_controller_v1_0.red;
     assign pixel_rgb[1] = hdmi_text_controller_v1_0.green;
     assign pixel_rgb[2] = hdmi_text_controller_v1_0.blue;
    
    // Pixel clock, hs, vs, and vde (!blank) - these come from your internal VGA module
     assign pixel_clk = hdmi_text_controller_v1_0.clk_25MHz;
     assign pixel_hs = hdmi_text_controller_v1_0.hsync;
     assign pixel_vs = hdmi_text_controller_v1_0.vsync;
     assign pixel_vde = hdmi_text_controller_v1_0.vde;
    
    // DrawX and DrawY - these come from your internal VGA module
     assign drawX = hdmi_text_controller_v1_0.drawX;
     assign drawY = hdmi_text_controller_v1_0.drawY;
   
    // BMP writing task, based off work from @BrianHGinc:
    // https://github.com/BrianHGinc/SystemVerilog-TestBench-BPM-picture-generator
    task save_bmp(string bmp_file_name);
        begin
        
            integer unsigned        fout_bmp_pointer, BMP_file_size,BMP_row_size,r;
            logic   unsigned [31:0] BMP_header[0:12];
        
                                      BMP_row_size  = 32'(BMP_WIDTH) & 32'hFFFC;  // When saving a bitmap, the row size/width must be
        if ((BMP_WIDTH & 32'd3) !=0)  BMP_row_size  = BMP_row_size + 4;           // padded to chunks of 4 bytes.
    
        fout_bmp_pointer= $fopen(bmp_file_name,"wb");
        if (fout_bmp_pointer==0) begin
            $display("Could not open file '%s' for writing",bmp_file_name);
            $stop;     
        end
        $display("Saving bitmap '%s'.",bmp_file_name);
       
        BMP_header[0:12] = '{BMP_file_size,0,0054,40,BMP_WIDTH,BMP_HEIGHT,{16'd24,16'd8},0,(BMP_row_size*BMP_HEIGHT*3),2835,2835,0,0};
        
        //Write header out      
        $fwrite(fout_bmp_pointer,"BM");
        for (int i =0 ; i <13 ; i++ ) $fwrite(fout_bmp_pointer,"%c%c%c%c",BMP_header[i][7 -:8],BMP_header[i][15 -:8],BMP_header[i][23 -:8],BMP_header[i][31 -:8]); // Better compatibility with Lattice Active_HDL.
        
        //Write image out (note that image is flipped in Y)
        for (int y=BMP_HEIGHT-1;y>=0;y--) begin
          for (int x=0;x<BMP_WIDTH;x++)
            $fwrite(fout_bmp_pointer,"%c%c%c",bitmap[x][y][23:16],bitmap[x][y][15:8],bitmap[x][y][7:0]) ;
        end
    
        $fclose(fout_bmp_pointer);
        end
    endtask
    
    // Always procedure to log RGB values into array to generate image
    always@(posedge pixel_clk)
        if (!arstn) begin
            for (j = 0; j < BMP_HEIGHT; j++)    //assign bitmap default to some light gray so we 
                for (i = 0; i < BMP_WIDTH; i++) //can tell the difference between drawn black
                    bitmap[i][j] <= 24'h0F0F0F; //and default color
        end
        else
            if (pixel_vde) //Only draw when not in the blanking interval
                bitmap[drawX][drawY] <= {pixel_rgb[0], 4'h0, pixel_rgb[1], 4'h0, pixel_rgb[2], 4'h00};
  
    // Provided AXI write task, follow this example for AXI read below
task axi_write_vram (
    input logic [11:0] addr, 
    input logic [6:0] code0, input logic [3:0] fgd_idx0, input logic [3:0] bkg_idx0, input logic iv0,
    input logic [6:0] code1, input logic [3:0] fgd_idx1, input logic [3:0] bkg_idx1, input logic iv1
);
    logic [31:0] data;
begin
    // Pack the data according to Table 7 format
    data = {iv1, code1, fgd_idx1, bkg_idx1, iv0, code0, fgd_idx0, bkg_idx0};
    
    $display("Writing data %h", data);
    
    // Perform AXI write with packed data
    #3 write_addr <= addr;        // Put write address on bus
    write_data <= data;           // Put packed data on bus
    write_addr_valid <= 1'b1;     // Indicate address is valid
    write_data_valid <= 1'b1;     // Indicate data is valid
    write_resp_ready <= 1'b1;     // Indicate ready for a response
    write_strb <= 4'hF;           // Writing all 4 bytes

    // Wait for slave ready signals or both signals and a positive edge clock
    wait(write_data_ready || write_addr_ready);
    @(posedge aclk);

    if(write_data_ready && write_addr_ready) begin
        write_addr_valid <= 0;
        write_data_valid <= 0;
    end else begin
        if(write_data_ready) begin
            write_data_valid <= 0;
            wait(write_addr_ready);
        end else if(write_addr_ready) begin
            write_addr_valid <= 0;
            wait(write_data_ready);
        end

        @(posedge aclk); // Complete second handshake
        write_addr_valid <= 0;
        write_data_valid <= 0;
    end

    // Deassert strobe and wait for valid response
    write_strb <= 4'h0;
    wait(write_resp_valid);
    @(posedge aclk);
    write_resp_ready <= 0;       // End of transaction
end
endtask

task axi_write_palette (
    input logic [31:0] addr,
    input logic [11:0] color1,   // First color (C1) in RGB format (12-bit)
    input logic [11:0] color2    // Second color (C2) in RGB format (12-bit)
);
    logic [31:0] data;
begin
    // Pack two colors into a single word (C1 in upper bits and C2 in lower bits)
    data = {6'b000000, color1[11:8], color1[7:4], color1[3:0], color2[11:8], color2[7:4], color2[3:0], 1'b0};
    
    #3 write_addr <= addr;              // Put address on bus (palette register address)
    write_data <= data;                 // Put packed colors on bus
    write_addr_valid <= 1'b1;           // Indicate address is valid
    write_data_valid <= 1'b1;           // Indicate data is valid
    write_resp_ready <= 1'b1;           // Indicate ready for response
    write_strb <= 4'hF;                 // Writing all bytes

    wait(write_data_ready || write_addr_ready);
    @(posedge aclk);

    if (write_data_ready && write_addr_ready) begin
        write_addr_valid <= 0;
        write_data_valid <= 0;
    end else begin
        if (write_data_ready) begin
            write_data_valid <= 0;
            wait(write_addr_ready);
        end else if (write_addr_ready) begin
            write_addr_valid <= 0;
            wait(write_data_ready);
        end

        @(posedge aclk);          // Complete second handshake
        write_addr_valid <= 0;
        write_data_valid <= 0;
    end

    wait(write_resp_valid);
    
    @(posedge aclk);    
    write_resp_ready <= 0;              // End of transaction   
end 
endtask

    
    //Fill in this task to perform an AXI read, similar to the provided example
    //of the AXI write above, follow the waveforms provided into the I.AMM manual
    //Note the read handshake process is simpler than the write
    task axi_read (input logic [31:0] addr, output logic [31:0] data);
        begin
            // Step 1: Initiate Read Address Phase
                read_addr <= addr;       // Set read address
                read_addr_valid <= 1'b1; // Indicate that address is valid
                
                // Wait for slave to assert ARREADY signal
                wait (read_addr_ready);
                
                // Step 2: Complete Address Handshake
                @(posedge aclk);         // Wait for clock edge
                read_addr_valid <= 1'b0; // Deassert ARVALID after handshake
                
                // Assert RREADY early, indicating readiness to accept data 
                read_data_ready <= 1'b1;
                
                // Step 3: Wait for Data Phase
                wait (read_data_valid);  // Wait for RVALID from slave
            
                // Step 4: Capture Data and Complete Data Handshake
                @(posedge aclk);         // Wait for clock edge
                data <= read_data;       // Capture data from RDATA
                
            
                @(posedge aclk);         // Wait for clock edge
                read_data_ready <= 1'b0; // Deassert RREADY after handshake
            
        end
    endtask;
  
  
    // Initial block for test vectors begins below
    initial begin: TEST_VECTORS
        arstn = 0; //reset IP
        repeat (4) @(posedge aclk);
        arstn <= 1;
        
        //remember AXI addresses are BYTE addresses!
  // Command 1: Black and Blue
// Write Blue and Green to the palette
repeat (4) @(posedge aclk) axi_write_palette(32'h2000, 12'h00F /* Blue */, 12'h00F /* Green */);

// Command 2: Green and Cyan
repeat (4) @(posedge aclk) axi_write_palette(32'h2004, 12'h0A0 /* Green */, 12'h0AA /* Cyan */);

// Command 3: Red and Magenta
repeat (4) @(posedge aclk) axi_write_palette(32'h2008, 12'hA00 /* Red */, 12'hA0A /* Magenta */);

// Command 4: Brown and Light Gray
repeat (4) @(posedge aclk) axi_write_palette(32'h200C, 12'hA50 /* Brown */, 12'hAAA /* Light Gray */);

// Command 5: Dark Gray and Light Blue
repeat (4) @(posedge aclk) axi_write_palette(32'h2010, 12'h555 /* Dark Gray */, 12'h55F /* Light Blue */);

// Command 6: Light Green and Light Cyan
repeat (4) @(posedge aclk) axi_write_palette(32'h2014, 12'h5F5 /* Light Green */, 12'h5FF /* Light Cyan */);

// Command 7: Light Red and Light Magenta
repeat (4) @(posedge aclk) axi_write_palette(32'h2018, 12'hF55 /* Light Red */, 12'hF5F /* Light Magenta */);

// Command 8: Yellow and White
repeat (4) @(posedge aclk) axi_write_palette(32'h201C, 12'hFF5 /* Yellow */, 12'hFFF /* White */);

            
            //Write into every one of the 600 VRAM registers, note that this is different than what the driver C code does
            //because the testbench axi_write task only generates aligned (full 32-bit) AXI writes (e.g. write_strb is always F)
            //The C code on the MicroBlaze expects to be able to do byte and halfword (16-bit) writes, therefore if the
            //simulation works but the checksum does not pass in the hardware, check handling of write_strb. 
    //        for(i=0; i < 1200; i++) begin 
    //		  repeat (4) @(posedge aclk) axi_write(4*i, i);
    //        end
            
            //The following is the readback routine. It tests that your AXI IP is capable of reading back all 601
            //VRAM registers via AXI (once you've properly filled in axi_read as above). Note that the verification
            //of the readback results is automatic, it will throw an assertion if the readback result is not as expected        
            ////////////////////////////////////////////
       /// Test Writing and Reading VRAM Entries //
       ////////////////////////////////////////////

       // Write "ansht2" in blue (foreground index = 1)
axi_write_vram(12'h000, /* ASCII 'a' */ 7'h61, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1,
                       /* ASCII 'n' */ 7'h6E, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1);

axi_write_vram(12'h004, /* ASCII 's' */ 7'h73, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1,
                       /* ASCII 'h' */ 7'h68, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1);

axi_write_vram(12'h008, /* ASCII 't' */ 7'h74, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1,
                       /* ASCII '2' */ 7'h32, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd1, /* IV */ 1'b1);
                       

               
// Write "completed" in red (foreground index = 3)
axi_write_vram(12'h012, /* ASCII 'c' */ 7'h63, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd0, /* IV */ 1'b1,
                       /* ASCII 'o' */ 7'h6F, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd0, /* IV */ 1'b1);

axi_write_vram(12'h016, /* ASCII 'm' */ 7'h6D, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd0, /* IV */ 1'b1,
                       /* ASCII 'p' */ 7'h70, /* FGD_IDX */ 4'd3, /* BKG_IDX */ 4'd0, /* IV */ 1'b1);

axi_write_vram(12'h01A, /* ASCII 'l' */ 7'h6C ,/*FGD_IDX*/4'd3 ,/*BKG*/4'd0 ,/*IV*/'b1,
                        /*ASCII 'e'*/7'h65 ,/*FGD*/4'd3 ,/*BKG*/'b0 ,/*IV*/'b1);

axi_write_vram(12'h01F ,/*ASCII 't'*/7'h74 ,/*FGD*/4'd3 ,/*BKG*/0 ,/*IV*/'b1,
                        /*ASCII 'e'*/7'h65 ,/*FGD*/4'd3 ,/*BKG*/0 ,/*IV*/'b1);

axi_write_vram(12'h023 ,/*ASCII 'd'*/7'h64 ,/*FGD*/4'd3 ,/*BKG*/0 ,/*IV*/'b1,
                        /*ASCII null (end)*/7'h00 ,/*FGD*/4'd3 ,/*BKG*/0 ,/*IV*/'b1);

// Write "ECE 385!" in green (foreground index = 2)
axi_write_vram(12'h027, /* ASCII 'E' */ 7'h45, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1,
                       /* ASCII 'C' */ 7'h43, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1);

axi_write_vram(12'h02B, /* ASCII 'E' */ 7'h45, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1,
                       /* ASCII '3' */ 7'h33, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1);

axi_write_vram(12'h02F, /* ASCII '8' */ 7'h38, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1,
                       /* ASCII '5'*/7'h35 ,/*FGD_IDX*/4'd2 ,/*BKG*/4'd0 ,/*IV*/'b01);

 axi_write_vram(12'h03C, /* ASCII '!' */ 7'h21, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1, /* ASCII '!' */ 7'h00, /* FGD_IDX */ 4'd2, /* BKG_IDX */ 4'd0, /* IV */ 1'b1);
    
       ////////////////////////////////////////
       /// Test Reading Back VRAM Entries   ///
       ////////////////////////////////////////

       for(i= 'd00;i<600;i++)begin 
            repeat(4)@(posedge aclk);
            axi_read(4*i,tb_read);

            axi_read_assert : assert(tb_read == {i+65,i%'d16,(i+8)%'d16,'b00,i+97,(i+8)%'d16,i%'d16,'b01})
                else $error("Mismatch at address %x. Expected:%h Actual:%h", i*4,{i+65,i%'d16,(i+8)%'d16,'b00,i+97,(i+8)%'d16,i%'d16,'b01},tb_read);
       end 
        
            
        repeat (4) @(posedge aclk) axi_read(600*4, tb_read);
        $info ("Read back of control register: %x", tb_read);
        
        //Make sure you've set the simulation settings to run to 'all', rather than the 1000ns default
		
		//Simulate until VS goes low (indicating a new frame) and write the results
		`ifdef SIM_VIDEO
		wait (drawY > 'h010);
		save_bmp ("lab7_1_sim.bmp");
		`endif
		$finish();
	end
    
endmodule	

	